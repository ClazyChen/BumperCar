﻿------------------------------------------
 -- 主程序
 -- 创建日期：2018-5-15
 -- 负责人：--
 -- 信号说明：
 --
------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity BumperCar is
	port(
		
